hjghjghujgvlgyv
